module nand5_delay (
    input  logic in1,
    input  logic in2,
    input  logic in3,
    input  logic in4,
    input  logic in5,
    output logic out
);
  //TODO: Complete the code
endmodule
