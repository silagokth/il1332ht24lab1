module propagate_logic (
    input  logic a,
    input  logic b,
    output logic p
);
  // TODO: Complete the code
endmodule
