module generate_logic (
    input  logic a,
    input  logic b,
    output logic g
);
  // TODO: Complete the code
endmodule
