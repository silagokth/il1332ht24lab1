module sum_logic (
    input  logic a,
    input  logic b,
    output logic carry_in,
    output logic sum
);
  //TODO: Complete the code
endmodule
